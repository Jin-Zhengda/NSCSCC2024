module cpu_axi (
    
);
    
endmodule