`timescale 1ns / 1ps
`include "core_defines.sv"
`include "csr_defines.sv"

module main_ex
    import pipeline_types::*;
(
    input dispatch_ex_t ex_i,

    // push forward
    input csr_push_forward_t mem_csr_pf,
    input csr_push_forward_t wb_csr_pf,

    // from csr
    input logic LLbit,

    // with dcache
    mem_dcache dcache_master,

    // with div
    ex_div div_master,

    // to bpu
    output branch_update update_info,

    // to ctrl
    output logic pause_alu,
    output logic branch_flush,

    // to dispatch
    output alu_op_t pre_ex_aluop,

    // to cache
    output cache_inst_t cache_inst,

    // to mem
    output ex_mem_t ex_o
);

    assign ex_o.pc = ex_i.pc;
    assign ex_o.inst = ex_i.inst;
    assign ex_o.inst_valid = ex_i.inst_valid;
    assign ex_o.is_privilege = ex_i.is_privilege;
    assign ex_o.aluop = ex_i.aluop;

    logic ex_is_exception;
    exception_cause_t ex_exception_cause;

    assign ex_o.is_exception = {ex_i.is_exception[5: 2], ex_is_exception, ex_i.is_exception[0]};
    assign ex_o.exception_cause = {ex_i.exception_cause[5: 2], ex_exception_cause, ex_i.exception_cause[0]};

    // regular alu
    bus32_t regular_alu_res;

    regular_alu u_regular_alu(
        .aluop(ex_i.aluop),
        .alusel(ex_i.alusel),

        .reg1(ex_i.reg1),
        .reg2(ex_i.reg2),

        .result(regular_alu_res)
    );
   
    // div alu
    logic pause_ex_div;
    logic start_div;
    logic op;
    logic done;

    bus32_t remainder;
    bus32_t quotient;

    assign start_div = (ex_i.aluop == `ALU_DIVW || ex_i.aluop == `ALU_MODW || ex_i.aluop == `ALU_DIVWU 
                        || ex_i.aluop == `ALU_MODWU) && !done;
    assign op = (ex_i.aluop == `ALU_DIVW || ex_i.aluop == `ALU_MODW);
    assign pause_ex_div = start_div;

    div_alu u_div_alu(
        .clk,
        .rst,

        .op,
        .dividend(ex_i.reg1),
        .divisor(ex_i.reg2),
        .start(start_div),

        .quotient_out(quotient),
        .remainder_out(remainder),
        .done
    );

    // branch alu
    bus32_t branch_alu_res;

    branch_alu u_branch_alu(
        .pc(ex_i.pc),
        .inst(ex_i.inst),
        .aluop(ex_i.aluop),

        .reg1(ex_i.reg1),
        .reg2(ex_i.reg2),

        .pre_is_branch_taken(ex_i.pre_is_branch_taken),
        .pre_branch_addr(ex_i.pre_branch_addr),

        .update_info(update_info),
        .branch_flush(branch_flush),
        .branch_alu_res(branch_alu_res)
    );

    // load store alu
    bus32_t load_store_alu_res;
    assign load_store_alu_res = (ex_i.aluop == `ALU_SCW)? {31'b0, LLbit}: 32'b0;

    logic is_mem;
    assign is_mem = ex_i.aluop == `ALU_LDB || ex_i.aluop == `ALU_LDBU || ex_i.aluop == `ALU_LDH 
                        || ex_i.aluop == `ALU_LDH || ex_i.aluop == `ALU_LDW || ex_i.aluop == `ALU_LLW
                        || ex_i.aluop == `ALU_PRELD || ex_i.aluop == `ALU_CACOP || ex_i.aluop == `ALU_STB
                        || ex_i.aluop == `ALU_STH || ex_i.aluop == `ALU_STW || ex_i.aluop == `ALU_SCW;

    logic pause_ex_mem;
    assign pause_ex_mem = is_mem && dcache_master.valid && !dcache_master.addr_ok;

    logic[11: 0] si12;
    logic[13: 9] si14;
    assign si12 = ex_i.inst[21: 10];
    assign si14 = ex_i.inst[14: 10];

    always_comb begin
        case (ex_i.aluop)
            `ALU_LDB, `ALU_LDBU, `ALU_LDH, `ALU_LDHU, `ALU_LDW, `ALU_LLW, `ALU_PRELD, `ALU_CACOP: begin
                ex_o.mem_addr = ex_i.reg1 + ex_i.reg2;
            end
            `ALU_STB, `ALU_STH, `ALU_STW: begin
                ex_o.mem_addr = ex_i.reg1 + {{20{si12[11]}}, si12};
            end
            `ALU_SCW: begin
                ex_o.mem_addr = ex_i.reg1 + {{16{si14[13]}}, si14, 2'b00};
            end
            default: begin
                ex_o.mem_addr = 32'b0;        
            end
        endcase
    end

    assign dcache_master.virtual_addr = ex_o.mem_addr;
    logic mem_is_valid;

    always_comb begin
        if (ex_o.is_exception == 6'b0) begin
            // if (ex_i.pc < 32'h1c000100) begin
            if (ex_i.pc < 32'h00000120) begin
                dcache_master.uncache_en = mem_is_valid;
                dcache_master.valid = 1'b0;
            end 
            else begin
                dcache_master.uncache_en = 1'b0;
                dcache_master.valid = mem_is_valid;
            end
        end
        else begin
            dcache_master.uncache_en = 1'b0;
            dcache_master.valid = 1'b0;
        end
    end

    always_comb begin: to_dcache
        case (ex_i.aluop) 
            `ALU_LDB, `ALU_LDBU: begin
                ex_is_exception = 1'b0;
                ex_exception_cause = 7'b0;
                dcache_master.op = 1'b0;
                mem_is_valid = 1'b1;
                dcache_master.wdata = 32'b0;
                dcache_master.wstrb = 4'b1111;
            end
            `ALU_LDH, `ALU_LDHU: begin
                ex_is_exception = ex_o.mem_addr[1: 0] == 2'b01 || ex_o.mem_addr[1: 0] == 2'b11;
                ex_exception_cause = (ex_o.mem_addr[1: 0] == 2'b01 || ex_o.mem_addr[1: 0] == 2'b11) ? `EXCEPTION_ALE : 7'b0;
                dcache_master.op = 1'b0;
                mem_is_valid = 1'b1;
                dcache_master.wdata = 32'b0;
                dcache_master.wstrb = 4'b1111;
            end
            `ALU_LDW, `ALU_LLW: begin
                ex_is_exception = ex_o.mem_addr[1: 0] == 2'b00;
                ex_exception_cause = (ex_o.mem_addr[1: 0] == 2'b00) ? 7'b0 : `EXCEPTION_ALE;
                dcache_master.op = 1'b0;
                mem_is_valid = 1'b1;
                dcache_master.wdata = 32'b0;
                dcache_master.wstrb = 4'b1111;
            end
            `ALU_STB: begin
                ex_is_exception = 1'b0;
                ex_exception_cause = 7'b0;
                dcache_master.op = 1'b1;
                dcache_master.wdata = {4{ex_i.reg2[7: 0]}};
                mem_is_valid = 1'b1;
                case (ex_o.mem_addr[1: 0])
                    2'b00: begin
                        dcache_master.wstrb = 4'b0001;
                    end 
                    2'b01: begin
                        dcache_master.wstrb = 4'b0010;
                    end
                    2'b10: begin
                        dcache_master.wstrb = 4'b0100;
                    end
                    2'b11: begin
                        dcache_master.wstrb = 4'b1000;
                    end
                    default: begin
                        dcache_master.wstrb = 4'b0000;                        
                    end
                endcase
            end
            `ALU_STH: begin
                dcache_master.op = 1'b1;
                dcache_master.wdata = {2{ex_i.reg2[15: 0]}};
                mem_is_valid = 1'b1;
                case (ex_o.mem_addr[1: 0])
                    2'b00: begin
                        dcache_master.wstrb = 4'b0011;
                        ex_is_exception = 1'b0;
                        ex_exception_cause = 7'b0;
                    end 
                    2'b10: begin
                        dcache_master.wstrb = 4'b1100;
                        ex_is_exception = 1'b0;
                        ex_exception_cause = 7'b0;
                    end
                    2'b01, 2'b11: begin
                        dcache_master.wstrb = 4'b0000;
                        ex_is_exception = 1'b1;
                        ex_exception_cause = `EXCEPTION_ALE;
                    end
                    default: begin
                        dcache_master.wstrb = 4'b0000;    
                        ex_is_exception = 1'b0;
                        ex_exception_cause = 7'b0;                    
                    end
                endcase
            end
            `ALU_STW: begin
                ex_is_exception = (ex_o.mem_addr[1: 0] == 2'b00) ? 1'b0 : 1'b1;
                ex_exception_cause = (ex_o.mem_addr[1: 0] == 2'b00) ? 7'b0 : `EXCEPTION_ALE;
                dcache_master.op = 1'b1;
                dcache_master.wdata = ex_i.reg2;
                mem_is_valid = 1'b1;
                dcache_master.wstrb = 4'b1111;
            end
            `ALU_SCW: begin
                ex_is_exception = (ex_o.mem_addr[1: 0] == 2'b00) ? 1'b0 : 1'b1;
                ex_exception_cause = (ex_o.mem_addr[1: 0] == 2'b00) ? 7'b0 : `EXCEPTION_ALE;
                if (LLbit) begin
                    dcache_master.op = 1'b1;
                    dcache_master.wdata = ex_i.reg2;
                    mem_is_valid = 1'b1;
                    dcache_master.wstrb = 4'b1111;
                end
                else begin
                    dcache_master.op = 1'b0;
                    dcache_master.wdata = 32'b0;
                    mem_is_valid = 1'b0;
                    dcache_master.wstrb = 4'b1111;
                end
            end
            default: begin
                mem_is_valid = 1'b0;
                dcache_master.wdata = 32'b0;
                dcache_master.op = 1'b0;
                dcache_master.wstrb = 4'b1111;
                ex_is_exception = 1'b0;
                ex_exception_cause = 7'b0;
            end
        endcase
    end

    always_comb begin
        if (ex_i.aluop == `ALU_LLW) begin
            ex_o.csr_write_en = 1'b1;
            ex_o.csr_addr = `CSR_LLBCTL;
            ex_o.csr_write_data = 32'b1;
            ex_o.is_llw_scw = 1'b1;
        end
        else if (ex_i.aluop == `ALU_SCW && LLbit) begin
            ex_o.csr_write_en = 1'b1;
            ex_o.csr_addr = `CSR_LLBCTL;
            ex_o.csr_write_data = 1'b0;
            ex_o.is_llw_scw = 1'b1;
        end
        else begin
            ex_o.csr_write_en = ex_i.csr_write_en;
            ex_o.csr_addr = ex_i.csr_addr;
            ex_o.csr_write_data = ex_i.reg1;
            ex_o.is_llw_scw = 1'b0;
        end
    end

    always_comb begin
        case (ex_i.aluop)
            `ALU_PRELD: begin
                cache_inst.is_cacop = 1'b0;
                cache_inst.cacop_code = 5'b0;
                cache_inst.is_preld = 1'b1;
                cache_inst.addr = ex_o.mem_addr;  
            end
            `ALU_CACOP: begin
                cache_inst.is_cacop = 1'b1;
                cache_inst.cacop_code = ex_i.cacop_code;
                cache_inst.is_preld = 1'b0;
                cache_inst.addr = ex_o.mem_addr;
            end
            default: begin
                cache_inst.is_cacop = 1'b0;
                cache_inst.cacop_code = 5'b0;
                cache_inst.is_preld = 1'b0;
                cache_inst.addr = 32'b0;
            end
        endcase
    end

    // csr alu
    bus32_t csr_alu_res;
    bus32_t csr_mask;


    // reg data 
    assign ex_o.reg_write_en = ex_i.reg_write_en;
    assign ex_o.reg_write_addr = ex_i.reg_write_addr;
    
    always_comb begin: reg_write
        case (ex_i.alusel)
            `ALU_SEL_LOGIC, `ALU_SEL_SHIFT,`ALU_SEL_ARITHMETIC: begin
                ex_o.reg_write_data = regular_alu_res;
            end
            `ALU_SEL_JUMP_BRANCH: begin
                ex_o.reg_write_data = branch_alu_res;
            end
            `ALU_SEL_LOAD_STORE: begin
                ex_o.reg_write_data = load_store_alu_res;
            end
            default: begin
                ex_o.reg_write_data = LLbit;
            end
        endcase
    end

    assign pause_alu = pause_ex_div || pause_ex_mem;

endmodule