`timescale 1ns / 1ps

module backend_top 
    import pipeline_types::*;
(
    input logic clk,
    input logic rst,

    input bus32_t pc,
    input logic inst,
    input logic pre_is_branch,
    input logic pre_is_branch_taken,
    input bus32_t pre_branch_addr,
    input logic [5:0] is_exception,
    input logic [5:0][EXC_CAUSE_WIDTH - 1:0] exception_cause,

    mem_dcache dcache_master,
    output cache_inst_t cache_inst
);

    // reg
    dispatch_regfile dispatch_regfile_io();

    // 
    
endmodule