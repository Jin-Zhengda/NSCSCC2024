module ram (
    
);
    
endmodule