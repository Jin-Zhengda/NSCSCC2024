`ifndef CSR_DEFINES_SV
`define CSR_DEFINES_SV

// CSR addresses
`define CSR_CRMD 14'b00000000000000
`define CSR_PRMD 14'b00000000000001
`define CSR_EUEN 14'b00000000000010
`define CSR_ECFG 14'b00000000000100
`define CSR_ESTAT 14'b00000000000101
`define CSR_ERA 14'b00000000000110
`define CSR_BADV 14'b00000000000111
`define CSR_EENTRY 14'b00000000001100
`define CSR_TLBIDX 14'b00000000010000
`define CSR_TLBHI 14'b00000000010001
`define CSR_TLBLO0 14'b00000000010010
`define CSR_TLBLO1 14'b00000000010011
`define CSR_ASID 14'b00000000011000
`define CSR_PGDL 14'b00000000011001
`define CSR_PGDH 14'b00000000011010
`define CSR_PGD 14'b00000000011011
`define CSR_CPUID 14'b00000000100000
`define CSR_SAVE0 14'b00000000110000
`define CSR_SAVE1 14'b00000000110001
`define CSR_SAVE2 14'b00000000110010
`define CSR_SAVE3 14'b00000000110011
`define CSR_TID 14'b00000001000000
`define CSR_TCFG 14'b00000001000001
`define CSR_TVAL 14'b00000001000010
`define CSR_TICLR 14'b00000001000100
`define CSR_LLBCTL 14'b00000001100000
`define CSR_TLBRENTRY 14'b00000010001000
`define CSR_CTAG 14'b00000010011000
`define CSR_DMW0 14'b00000110000000
`define CSR_DMW1 14'b00000110000001

// Exceptions
`define EXCEPTION_INT 7'b0000000
`define EXCEPTION_PIL 7'b0000010
`define EXCEPTION_PIS 7'b0000100
`define EXCEPTION_PIF 7'b0000110
`define EXCEPTION_PME 7'b0001000
`define EXCEPTION_PPI 7'b0001110
`define EXCEPTION_ADEF 7'b0010000
`define EXCEPTION_ADEM  7'b0010001
`define EXCEPTION_ALE 7'b0010010
`define EXCEPTION_SYS 7'b0010110
`define EXCEPTION_BRK 7'b0011000
`define EXCEPTION_INE 7'b0011010
`define EXCEPTION_IPE 7'b0011100
`define EXCEPTION_FPD 7'b0011110
`define EXCEPTION_FPE 7'b0100100
`define EXCEPTION_TLBR 7'b1111110
`define EXCEPTION_NOP 7'b1111111

`endif