module cpu_top (
 
);